module fetch_tb();
/*
	logic PCSrc_F,clk,reset;
	logic [63:0] PCBranch_F,imem_addr_F
	
	fetch dut (PCSrc_F,clk,reset,PCBranch_F,imem_addr_F);

	always 
		begin
			5# clk = ~clk;
		end 
		
	initial
		begin
			reset = 1; #5;
			clk = 0; 
		end 
*/
endmodule 
